module ramWhithClock;

endmodule