module muxForM3AndM4Output(selectRegister,r0,r1,r2,r3,r4,r5,r6,r7)
endmodule
